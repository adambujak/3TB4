module lab1part1 ( input a, output b );
	
endmodule
