//D flip flop
module dff (input d,clk, output reg q, output q_b);
	always @(posedge clk)
	begin
		q<=d;
	end
	assign q_b = ~q;
endmodule

//D latch
module dlatch(data, en, q);
	output q;
	reg q; 
	always @(en or data)
	begin
		if (en)
			q <= data;
	end
endmodule

//4-1 MUX
module mux_4to1_case (input a, b, c, input [1:0] sel, output reg out); 
	always @ (*)
	begin
		case (sel)
		2'b00 : out <= a;
		2'b01 : out <= b;
		2'b10 : out <= c;
		2'b11 : out <= d;
		endcase
	end
endmodule

//4-bit counter
module counter(input clk, input rst, output reg[3:0] out);
	always @ (posedge clk)
	begin
		if(!rst)
			out <= 0;
		else
			out <= out + 1;
	end
endmodule
